library IEEE; 
use IEEE.STD_LOGIC_1164.ALL; 

ENTITY half_adder_e IS  --- Half Adder 
PORT(
a,b:in std_logic; 
s,c :out std_logic
); 
END half_adder_e; 
